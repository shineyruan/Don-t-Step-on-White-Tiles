///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: <Name>
//
// File: write_pos.v
// File history:
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//      <Revision number>: <Date>: <Comments>
//
// Description: 
//
// <Description here>
//
// Targeted device: <Family::SmartFusion> <Die::A2F200M3F> <Package::484 FBGA>
// Author: <Name>
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

//`timescale <time_units> / <precision>

module write_pos( port1, port2, port3, port4 );
input port1, port2;
output port3;
inout port4;

//<statements>

endmodule

