// Actel Corporation Proprietary and Confidential
// Copyright 2010 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
// Revision Information:
// 05Feb10              Production Release Version 3.0
// SVN Revision Information:
// SVN $Revision: 24054 $
// SVN $Date: 2014-12-08 10:43:40 +0000 (Mon, 08 Dec 2014) $
`timescale 1ns/1ps
module
CAPB3II
(
input
[
16
:
0
]
CAPB3lI,
input
[
31
:
0
]
PRDATAS0,
input
[
31
:
0
]
PRDATAS1,
input
[
31
:
0
]
PRDATAS2,
input
[
31
:
0
]
PRDATAS3,
input
[
31
:
0
]
PRDATAS4,
input
[
31
:
0
]
PRDATAS5,
input
[
31
:
0
]
PRDATAS6,
input
[
31
:
0
]
PRDATAS7,
input
[
31
:
0
]
PRDATAS8,
input
[
31
:
0
]
PRDATAS9,
input
[
31
:
0
]
PRDATAS10,
input
[
31
:
0
]
PRDATAS11,
input
[
31
:
0
]
PRDATAS12,
input
[
31
:
0
]
PRDATAS13,
input
[
31
:
0
]
PRDATAS14,
input
[
31
:
0
]
PRDATAS15,
input
[
31
:
0
]
PRDATAS16,
input
[
16
:
0
]
CAPB3Ol,
input
[
16
:
0
]
CAPB3Il,
output
wire
PREADY,
output
wire
PSLVERR,
output
wire
[
31
:
0
]
PRDATA
)
;
localparam
[
4
:
0
]
CAPB3ll
=
5
'b
00000
;
localparam
[
4
:
0
]
CAPB3O0
=
5
'b
00001
;
localparam
[
4
:
0
]
CAPB3I0
=
5
'b
00010
;
localparam
[
4
:
0
]
CAPB3l0
=
5
'b
00011
;
localparam
[
4
:
0
]
CAPB3O1
=
5
'b
00100
;
localparam
[
4
:
0
]
CAPB3I1
=
5
'b
00101
;
localparam
[
4
:
0
]
CAPB3l1
=
5
'b
00110
;
localparam
[
4
:
0
]
CAPB3OOI
=
5
'b
00111
;
localparam
[
4
:
0
]
CAPB3IOI
=
5
'b
01000
;
localparam
[
4
:
0
]
CAPB3lOI
=
5
'b
01001
;
localparam
[
4
:
0
]
CAPB3OII
=
5
'b
01010
;
localparam
[
4
:
0
]
CAPB3III
=
5
'b
01011
;
localparam
[
4
:
0
]
CAPB3lII
=
5
'b
01100
;
localparam
[
4
:
0
]
CAPB3OlI
=
5
'b
01101
;
localparam
[
4
:
0
]
CAPB3IlI
=
5
'b
01110
;
localparam
[
4
:
0
]
CAPB3llI
=
5
'b
01111
;
localparam
[
4
:
0
]
CAPB3O0I
=
5
'b
10000
;
reg
CAPB3I0I
;
reg
CAPB3l0I
;
reg
[
31
:
0
]
CAPB3O1I
;
wire
[
4
:
0
]
CAPB3I1I
;
wire
[
31
:
0
]
CAPB3l1I
;
assign
CAPB3l1I
=
32
'b
0
;
assign
CAPB3I1I
[
4
]
=
CAPB3lI
[
16
]
;
assign
CAPB3I1I
[
3
]
=
CAPB3lI
[
15
]
|
CAPB3lI
[
14
]
|
CAPB3lI
[
13
]
|
CAPB3lI
[
12
]
|
CAPB3lI
[
11
]
|
CAPB3lI
[
10
]
|
CAPB3lI
[
9
]
|
CAPB3lI
[
8
]
;
assign
CAPB3I1I
[
2
]
=
CAPB3lI
[
15
]
|
CAPB3lI
[
14
]
|
CAPB3lI
[
13
]
|
CAPB3lI
[
12
]
|
CAPB3lI
[
7
]
|
CAPB3lI
[
6
]
|
CAPB3lI
[
5
]
|
CAPB3lI
[
4
]
;
assign
CAPB3I1I
[
1
]
=
CAPB3lI
[
15
]
|
CAPB3lI
[
14
]
|
CAPB3lI
[
11
]
|
CAPB3lI
[
10
]
|
CAPB3lI
[
7
]
|
CAPB3lI
[
6
]
|
CAPB3lI
[
3
]
|
CAPB3lI
[
2
]
;
assign
CAPB3I1I
[
0
]
=
CAPB3lI
[
15
]
|
CAPB3lI
[
13
]
|
CAPB3lI
[
11
]
|
CAPB3lI
[
9
]
|
CAPB3lI
[
7
]
|
CAPB3lI
[
5
]
|
CAPB3lI
[
3
]
|
CAPB3lI
[
1
]
;
always
@
(
*
)
begin
case
(
CAPB3I1I
)
CAPB3ll
:
if
(
CAPB3lI
[
0
]
)
CAPB3O1I
[
31
:
0
]
=
PRDATAS0
[
31
:
0
]
;
else
CAPB3O1I
[
31
:
0
]
=
CAPB3l1I
[
31
:
0
]
;
CAPB3O0
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS1
[
31
:
0
]
;
CAPB3I0
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS2
[
31
:
0
]
;
CAPB3l0
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS3
[
31
:
0
]
;
CAPB3O1
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS4
[
31
:
0
]
;
CAPB3I1
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS5
[
31
:
0
]
;
CAPB3l1
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS6
[
31
:
0
]
;
CAPB3OOI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS7
[
31
:
0
]
;
CAPB3IOI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS8
[
31
:
0
]
;
CAPB3lOI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS9
[
31
:
0
]
;
CAPB3OII
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS10
[
31
:
0
]
;
CAPB3III
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS11
[
31
:
0
]
;
CAPB3lII
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS12
[
31
:
0
]
;
CAPB3OlI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS13
[
31
:
0
]
;
CAPB3IlI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS14
[
31
:
0
]
;
CAPB3llI
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS15
[
31
:
0
]
;
CAPB3O0I
:
CAPB3O1I
[
31
:
0
]
=
PRDATAS16
[
31
:
0
]
;
default
:
CAPB3O1I
[
31
:
0
]
=
CAPB3l1I
[
31
:
0
]
;
endcase
end
always
@
(
*
)
begin
case
(
CAPB3I1I
)
CAPB3ll
:
if
(
CAPB3lI
[
0
]
)
CAPB3I0I
=
CAPB3Ol
[
0
]
;
else
CAPB3I0I
=
1
'b
1
;
CAPB3O0
:
CAPB3I0I
=
CAPB3Ol
[
1
]
;
CAPB3I0
:
CAPB3I0I
=
CAPB3Ol
[
2
]
;
CAPB3l0
:
CAPB3I0I
=
CAPB3Ol
[
3
]
;
CAPB3O1
:
CAPB3I0I
=
CAPB3Ol
[
4
]
;
CAPB3I1
:
CAPB3I0I
=
CAPB3Ol
[
5
]
;
CAPB3l1
:
CAPB3I0I
=
CAPB3Ol
[
6
]
;
CAPB3OOI
:
CAPB3I0I
=
CAPB3Ol
[
7
]
;
CAPB3IOI
:
CAPB3I0I
=
CAPB3Ol
[
8
]
;
CAPB3lOI
:
CAPB3I0I
=
CAPB3Ol
[
9
]
;
CAPB3OII
:
CAPB3I0I
=
CAPB3Ol
[
10
]
;
CAPB3III
:
CAPB3I0I
=
CAPB3Ol
[
11
]
;
CAPB3lII
:
CAPB3I0I
=
CAPB3Ol
[
12
]
;
CAPB3OlI
:
CAPB3I0I
=
CAPB3Ol
[
13
]
;
CAPB3IlI
:
CAPB3I0I
=
CAPB3Ol
[
14
]
;
CAPB3llI
:
CAPB3I0I
=
CAPB3Ol
[
15
]
;
CAPB3O0I
:
CAPB3I0I
=
CAPB3Ol
[
16
]
;
default
:
CAPB3I0I
=
1
'b
1
;
endcase
end
always
@
(
*
)
begin
case
(
CAPB3I1I
)
CAPB3ll
:
if
(
CAPB3lI
[
0
]
)
CAPB3l0I
=
CAPB3Il
[
0
]
;
else
CAPB3l0I
=
1
'b
0
;
CAPB3O0
:
CAPB3l0I
=
CAPB3Il
[
1
]
;
CAPB3I0
:
CAPB3l0I
=
CAPB3Il
[
2
]
;
CAPB3l0
:
CAPB3l0I
=
CAPB3Il
[
3
]
;
CAPB3O1
:
CAPB3l0I
=
CAPB3Il
[
4
]
;
CAPB3I1
:
CAPB3l0I
=
CAPB3Il
[
5
]
;
CAPB3l1
:
CAPB3l0I
=
CAPB3Il
[
6
]
;
CAPB3OOI
:
CAPB3l0I
=
CAPB3Il
[
7
]
;
CAPB3IOI
:
CAPB3l0I
=
CAPB3Il
[
8
]
;
CAPB3lOI
:
CAPB3l0I
=
CAPB3Il
[
9
]
;
CAPB3OII
:
CAPB3l0I
=
CAPB3Il
[
10
]
;
CAPB3III
:
CAPB3l0I
=
CAPB3Il
[
11
]
;
CAPB3lII
:
CAPB3l0I
=
CAPB3Il
[
12
]
;
CAPB3OlI
:
CAPB3l0I
=
CAPB3Il
[
13
]
;
CAPB3IlI
:
CAPB3l0I
=
CAPB3Il
[
14
]
;
CAPB3llI
:
CAPB3l0I
=
CAPB3Il
[
15
]
;
CAPB3O0I
:
CAPB3l0I
=
CAPB3Il
[
16
]
;
default
:
CAPB3l0I
=
1
'b
0
;
endcase
end
assign
PREADY
=
CAPB3I0I
;
assign
PSLVERR
=
CAPB3l0I
;
assign
PRDATA
=
CAPB3O1I
[
31
:
0
]
;
endmodule
